-- touch contoller code


